library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

package constants is
	constant Nb : integer := 14;
	constant N : integer := 1;
 --  constant a1 : std_logic_vector (Nb-1 downto 0)  := "11101011101110"; --"00010100010010"; -- (= 1298)
--	constant b1 : std_logic_vector (Nb-1 downto 0) := "00110101110111"; -- (= 3447)
--	constant b0 : std_logic_vector (Nb-1 downto 0) := "00110101110111"; -- (= 3447)
--	constant a1b0 : std_logic_vector (23 downto 0) := "101110111011101010100010";--"010001000100010101011110"; -- (= 4474206) -> (-a1 * b0)
--	constant a1b1 : std_logic_vector (23 downto 0) := "101110111011101010100010"; --"010001000100010101011110"; -- (= 4474206) -> (-a1 * b1)

end constants;
