library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

package constants is
	constant Nb : integer := 14;
	constant N : integer := 1;
 --   constant a1 : signed (Nb-1 downto 0) :="11101011101110"; -- "111010"; --"11101011101110";
--	constant b1 : signed (Nb-1 downto 0) := "00110101110111"; -- "001101"; --"00110101110111";
--	constant b0 : signed (Nb-1 downto 0) :="00110101110111"; -- "001101"; --"00110101110111";
end constants;
